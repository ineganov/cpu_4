module testbench;
//====================================================================// 
logic       CLK, RESET;
logic [7:0] LEDS;
if_io IO();
//====================================================================// 
always
  begin
  CLK = ~CLK;
  #10ns;
  end 
//====================================================================// 
initial
  begin
  CLK = 0;
  RESET = 1;

  repeat(2)
    @(posedge CLK) #10;
  RESET = 0; 

  end
//====================================================================// 

mcpu   mcpu  (.CLK       ( CLK   ),
              .RESET     ( RESET ),
              .IO        ( IO    ));

ffd #(8) led_reg(CLK, RESET, IO.LEDS_WE, IO.LEDS_WD, LEDS);

//====================================================================// 
endmodule
